* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461702396344 1 2 4
** N=5 EP=3 IP=0 FDC=1
M0 2 5 1 4 nch L=2e-06 W=2.05e-06 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461702396342 1 2
** N=7 EP=2 IP=0 FDC=1
M0 2 5 1 6 pch L=5e-06 W=2e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461702396346 1 2 4
** N=5 EP=3 IP=0 FDC=1
M0 2 5 1 4 nch L=5e-06 W=2e-05 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461702396343 1
** N=7 EP=1 IP=0 FDC=1
M0 1 5 4 6 pch L=1e-06 W=2e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461702396349 1 2 4
** N=5 EP=3 IP=0 FDC=1
M0 2 5 1 4 nch L=2e-06 W=2e-05 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_4617023963410 1
** N=7 EP=1 IP=0 FDC=1
M0 1 5 4 6 pch L=1e-06 W=2.03e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461702396340 1 2 4
** N=5 EP=3 IP=0 FDC=1
M0 2 5 1 4 nch L=1e-06 W=2e-05 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461702396345 1
** N=7 EP=1 IP=0 FDC=1
M0 1 5 4 6 pch L=2e-06 W=2e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT comparator_rail2rail_input_external_current Gnd Out Ref In Vdd
** N=32 EP=5 IP=100 FDC=31
M0 Out 27 Gnd 30 nch L=5e-07 W=1e-06 $X=48070 $Y=20955 $D=28
M1 Out 28 3 31 pch L=5e-07 W=2e-06 $X=49280 $Y=25305 $D=62
X2 10 18 rppolywo l=3.831e-05 w=8e-07 $X=4870 $Y=2205 $D=215
X3 Gnd 9 30 nch_mac_CDNS_461702396344 $T=42090 19905 0 0 $X=41730 $Y=19545
X4 Gnd 9 30 nch_mac_CDNS_461702396344 $T=45080 19905 0 0 $X=44720 $Y=19545
X5 22 20 pch_mac_CDNS_461702396342 $T=36650 25305 0 0 $X=36200 $Y=24945
X6 22 25 pch_mac_CDNS_461702396342 $T=43050 25305 0 0 $X=42600 $Y=24945
X7 4 5 30 nch_mac_CDNS_461702396346 $T=29700 1955 0 0 $X=29340 $Y=1595
X8 4 6 30 nch_mac_CDNS_461702396346 $T=36100 1955 0 0 $X=35740 $Y=1595
X9 7 pch_mac_CDNS_461702396343 $T=14180 25305 0 0 $X=13730 $Y=24945
X10 8 pch_mac_CDNS_461702396343 $T=16410 25305 0 0 $X=15960 $Y=24945
X11 6 pch_mac_CDNS_461702396343 $T=27560 25305 0 0 $X=27110 $Y=24945
X12 6 pch_mac_CDNS_461702396343 $T=29790 25305 0 0 $X=29340 $Y=24945
X13 9 pch_mac_CDNS_461702396343 $T=32020 25305 0 0 $X=31570 $Y=24945
X14 9 pch_mac_CDNS_461702396343 $T=34250 25305 0 0 $X=33800 $Y=24945
X15 Gnd 10 30 nch_mac_CDNS_461702396349 $T=23310 1960 0 0 $X=22950 $Y=1600
X16 Gnd 4 30 nch_mac_CDNS_461702396349 $T=26300 1960 0 0 $X=25940 $Y=1600
X17 11 pch_mac_CDNS_4617023963410 $T=18640 25005 0 0 $X=18190 $Y=24645
X18 11 pch_mac_CDNS_4617023963410 $T=20870 25005 0 0 $X=20420 $Y=24645
X19 5 pch_mac_CDNS_4617023963410 $T=23100 25005 0 0 $X=22650 $Y=24645
X20 5 pch_mac_CDNS_4617023963410 $T=25330 25005 0 0 $X=24880 $Y=24645
X21 Gnd 12 30 nch_mac_CDNS_461702396340 $T=7390 1955 0 0 $X=7030 $Y=1595
X22 Gnd 13 30 nch_mac_CDNS_461702396340 $T=9380 1955 0 0 $X=9020 $Y=1595
X23 Gnd 11 30 nch_mac_CDNS_461702396340 $T=11370 1955 0 0 $X=11010 $Y=1595
X24 Gnd 11 30 nch_mac_CDNS_461702396340 $T=13360 1955 0 0 $X=13000 $Y=1595
X25 Gnd 5 30 nch_mac_CDNS_461702396340 $T=15350 1955 0 0 $X=14990 $Y=1595
X26 Gnd 5 30 nch_mac_CDNS_461702396340 $T=17340 1955 0 0 $X=16980 $Y=1595
X27 Gnd 14 30 nch_mac_CDNS_461702396340 $T=19330 1955 0 0 $X=18970 $Y=1595
X28 Gnd 15 30 nch_mac_CDNS_461702396340 $T=21320 1955 0 0 $X=20960 $Y=1595
X29 21 pch_mac_CDNS_461702396345 $T=7720 25305 0 0 $X=7270 $Y=24945
X30 22 pch_mac_CDNS_461702396345 $T=10950 25305 0 0 $X=10500 $Y=24945
.ENDS
***************************************
