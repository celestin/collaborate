* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461775348295
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461775348297
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_4617753482910
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461775348290
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461775348292
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_4617753482911
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461775348294
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461775348293
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461775348299
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT comparator_rail2rail_input_external_current Gnd Out Vdd In Ref
** N=14 EP=5 IP=100 FDC=31
M0 Out 7 Gnd Gnd nch L=5e-07 W=1e-06 AD=2.3e-13 AS=2.3e-13 PD=2.46e-06 PS=2.46e-06 NRD=0.23 NRS=0.23 sa=2.3e-07 sb=2.3e-07 sca=1.77318 scb=0.000164701 scc=8.24936e-08 $X=31695 $Y=22735 $D=28
M1 5 In 4 Gnd nch L=5e-07 W=2e-06 AD=4.6e-13 AS=4.6e-13 PD=4.46e-06 PS=4.46e-06 NRD=0.115 NRS=0.115 sa=2.3e-07 sb=2.3e-07 sca=0.322415 scb=9.93945e-08 scc=6.57835e-14 $X=29290 $Y=1960 $D=28
M2 6 Ref 4 Gnd nch L=5e-07 W=2e-06 AD=4.6e-13 AS=4.6e-13 PD=4.46e-06 PS=4.46e-06 NRD=0.115 NRS=0.115 sa=2.3e-07 sb=2.3e-07 sca=0.322415 scb=9.93945e-08 scc=6.57835e-14 $X=31280 $Y=1960 $D=28
M3 7 8 Gnd Gnd nch L=2e-06 W=5e-06 AD=1.15e-12 AS=1.15e-12 PD=1.046e-05 PS=1.046e-05 NRD=0.046 NRS=0.046 sa=2.3e-07 sb=2.3e-07 sca=0.0971429 scb=1.37713e-22 scc=1.31505e-44 $X=29290 $Y=5860 $D=28
M4 7 8 Gnd Gnd nch L=2e-06 W=5e-06 AD=1.15e-12 AS=1.15e-12 PD=1.046e-05 PS=1.046e-05 NRD=0.046 NRS=0.046 sa=2.3e-07 sb=2.3e-07 sca=0.205143 scb=1.0062e-07 scc=1.80543e-13 $X=29290 $Y=12195 $D=28
M5 8 8 Gnd Gnd nch L=2e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.109982 scb=9.93946e-09 scc=6.57835e-15 $X=23310 $Y=1960 $D=28
M6 4 8 Gnd Gnd nch L=2e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.183369 scb=1.20436e-05 scc=1.60631e-08 $X=26300 $Y=1960 $D=28
M7 9 9 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.115312 scb=1.0413e-08 scc=7.24424e-15 $X=7390 $Y=1955 $D=28
M8 9 9 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.115312 scb=1.0413e-08 scc=7.24424e-15 $X=9380 $Y=1955 $D=28
M9 6 9 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.115312 scb=1.0413e-08 scc=7.24424e-15 $X=11370 $Y=1955 $D=28
M10 6 9 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.115312 scb=1.0413e-08 scc=7.24424e-15 $X=13360 $Y=1955 $D=28
M11 5 10 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.115312 scb=1.0413e-08 scc=7.24424e-15 $X=15350 $Y=1955 $D=28
M12 5 10 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.116111 scb=1.0413e-08 scc=7.24424e-15 $X=17340 $Y=1955 $D=28
M13 10 10 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.116977 scb=1.0413e-08 scc=7.24424e-15 $X=19330 $Y=1955 $D=28
M14 10 10 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.116977 scb=1.0413e-08 scc=7.24424e-15 $X=21320 $Y=1955 $D=28
M15 Out 7 Vdd Vdd pch L=5e-07 W=2e-06 AD=4.6e-13 AS=6.4e-13 PD=4.46e-06 PS=4.64e-06 NRD=0.115 NRS=0.16 sa=5.6e-07 sb=2.3e-07 sca=7.43579 scb=0.00482332 scc=0.000171928 $X=33660 $Y=21735 $D=62
M16 5 5 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.516267 scb=0.00035457 scc=1.65744e-05 $X=14180 $Y=25305 $D=62
M17 6 6 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.517394 scb=0.00035457 scc=1.65744e-05 $X=29790 $Y=25305 $D=62
M18 7 6 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.584328 scb=0.00035457 scc=1.65744e-05 $X=32020 $Y=25305 $D=62
M19 7 6 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=2.0155 scb=0.000965487 scc=1.96597e-05 $X=34250 $Y=25305 $D=62
M20 9 In 12 Vdd pch L=5e-07 W=2e-06 AD=4.6e-13 AS=4.6e-13 PD=4.46e-06 PS=4.46e-06 NRD=0.115 NRS=0.115 sa=2.3e-07 sb=2.3e-07 sca=6.53892 scb=0.00475197 scc=0.000171914 $X=29335 $Y=18665 $D=62
M21 10 Ref 12 Vdd pch L=5e-07 W=2e-06 AD=4.6e-13 AS=4.6e-13 PD=4.46e-06 PS=4.46e-06 NRD=0.115 NRS=0.115 sa=2.3e-07 sb=2.3e-07 sca=4.97027 scb=0.00356126 scc=0.000165745 $X=31235 $Y=18665 $D=62
M22 5 5 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.516267 scb=0.00035457 scc=1.65744e-05 $X=16410 $Y=25305 $D=62
M23 6 6 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.516267 scb=0.00035457 scc=1.65744e-05 $X=27560 $Y=25305 $D=62
M24 6 5 Vdd Vdd pch L=1e-06 W=2.03e-05 AD=4.669e-12 AS=6.496e-12 PD=4.106e-05 PS=4.124e-05 NRD=0.01133 NRS=0.0157635 sa=5.6e-07 sb=2.3e-07 sca=0.512401 scb=0.000349472 scc=1.63295e-05 $X=18640 $Y=25005 $D=62
M25 6 5 Vdd Vdd pch L=1e-06 W=2.03e-05 AD=4.669e-12 AS=6.496e-12 PD=4.106e-05 PS=4.124e-05 NRD=0.01133 NRS=0.0157635 sa=5.6e-07 sb=2.3e-07 sca=0.509893 scb=0.00034933 scc=1.63295e-05 $X=20870 $Y=25005 $D=62
M26 5 6 Vdd Vdd pch L=1e-06 W=2.03e-05 AD=4.669e-12 AS=6.496e-12 PD=4.106e-05 PS=4.124e-05 NRD=0.01133 NRS=0.0157635 sa=5.6e-07 sb=2.3e-07 sca=0.509962 scb=0.00034933 scc=1.63295e-05 $X=23100 $Y=25005 $D=62
M27 5 6 Vdd Vdd pch L=1e-06 W=2.03e-05 AD=4.669e-12 AS=6.496e-12 PD=4.106e-05 PS=4.124e-05 NRD=0.01133 NRS=0.0157635 sa=5.6e-07 sb=2.3e-07 sca=0.515602 scb=0.000351738 scc=1.63416e-05 $X=25330 $Y=25005 $D=62
M28 11 11 Vdd Vdd pch L=2e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.939341 scb=0.000372598 scc=1.65779e-05 $X=7720 $Y=25305 $D=62
M29 12 11 Vdd Vdd pch L=2e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.519665 scb=0.00035457 scc=1.65744e-05 $X=10950 $Y=25305 $D=62
X30 8 11 rppolywo l=3.831e-05 w=8e-07 $X=4870 $Y=2205 $D=215
.ENDS
***************************************
