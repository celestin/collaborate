* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_4618498380410 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=1e-06 W=2e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_4618498380412 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 4 1 3 nch L=5e-07 W=2e-06 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_4618498380415 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 2 4 1 3 pch L=5e-07 W=2e-06 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461849838045 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=2e-06 W=5e-06 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461849838047 1 2
** N=3 EP=2 IP=0 FDC=1
M0 2 2 1 1 pch L=1e-06 W=2e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_4618498380416 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=2e-06 W=2e-05 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461849838049 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=1e-06 W=2.03e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461849838048 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=1e-06 W=2e-05 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_4618498380414 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=2e-06 W=2e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT comparator_rail2rail_input_external_current Gnd Out Vdd In Ref
** N=14 EP=5 IP=100 FDC=31
M0 Out 9 Gnd Gnd nch L=5e-07 W=1e-06 $X=31695 $Y=22735 $D=28
M1 Out 9 Vdd Vdd pch L=5e-07 W=2e-06 $X=33660 $Y=21735 $D=62
X2 10 13 rppolywo l=3.831e-05 w=8e-07 $X=4870 $Y=2205 $D=215
X3 Vdd 7 7 pch_mac_CDNS_4618498380410 $T=14180 25305 0 0 $X=13400 $Y=24945
X4 Vdd 8 8 pch_mac_CDNS_4618498380410 $T=29790 25305 0 0 $X=29010 $Y=24945
X5 Vdd 9 8 pch_mac_CDNS_4618498380410 $T=32020 25305 0 0 $X=31240 $Y=24945
X6 Vdd 9 8 pch_mac_CDNS_4618498380410 $T=34250 25305 0 0 $X=33470 $Y=24945
X7 6 7 Gnd In nch_mac_CDNS_4618498380412 $T=29290 1960 0 0 $X=28930 $Y=1600
X8 6 8 Gnd Ref nch_mac_CDNS_4618498380412 $T=31280 1960 0 0 $X=30920 $Y=1600
X9 14 11 Vdd In pch_mac_CDNS_4618498380415 $T=29335 18665 0 0 $X=28885 $Y=18145
X10 14 12 Vdd Ref pch_mac_CDNS_4618498380415 $T=31235 18665 0 0 $X=30785 $Y=18145
X11 Gnd 9 10 nch_mac_CDNS_461849838045 $T=29290 5860 0 0 $X=28930 $Y=5340
X12 Gnd 9 10 nch_mac_CDNS_461849838045 $T=29290 12195 0 0 $X=28930 $Y=11675
X13 Vdd 7 pch_mac_CDNS_461849838047 $T=16410 25305 0 0 $X=15630 $Y=24785
X14 Vdd 8 pch_mac_CDNS_461849838047 $T=27560 25305 0 0 $X=26780 $Y=24785
X15 Gnd 10 10 nch_mac_CDNS_4618498380416 $T=23310 1960 0 0 $X=22950 $Y=1600
X16 Gnd 6 10 nch_mac_CDNS_4618498380416 $T=26300 1960 0 0 $X=25940 $Y=1600
X17 Vdd 8 7 pch_mac_CDNS_461849838049 $T=18640 25005 0 0 $X=17860 $Y=24645
X18 Vdd 8 7 pch_mac_CDNS_461849838049 $T=20870 25005 0 0 $X=20090 $Y=24645
X19 Vdd 7 8 pch_mac_CDNS_461849838049 $T=23100 25005 0 0 $X=22320 $Y=24645
X20 Vdd 7 8 pch_mac_CDNS_461849838049 $T=25330 25005 0 0 $X=24550 $Y=24645
X21 Gnd 11 11 nch_mac_CDNS_461849838048 $T=7390 1955 0 0 $X=7030 $Y=1595
X22 Gnd 11 11 nch_mac_CDNS_461849838048 $T=9380 1955 0 0 $X=9020 $Y=1595
X23 Gnd 8 11 nch_mac_CDNS_461849838048 $T=11370 1955 0 0 $X=11010 $Y=1595
X24 Gnd 8 11 nch_mac_CDNS_461849838048 $T=13360 1955 0 0 $X=13000 $Y=1595
X25 Gnd 7 12 nch_mac_CDNS_461849838048 $T=15350 1955 0 0 $X=14990 $Y=1595
X26 Gnd 7 12 nch_mac_CDNS_461849838048 $T=17340 1955 0 0 $X=16980 $Y=1595
X27 Gnd 12 12 nch_mac_CDNS_461849838048 $T=19330 1955 0 0 $X=18970 $Y=1595
X28 Gnd 12 12 nch_mac_CDNS_461849838048 $T=21320 1955 0 0 $X=20960 $Y=1595
X29 Vdd 13 13 pch_mac_CDNS_4618498380414 $T=7720 25305 0 0 $X=6940 $Y=24945
X30 Vdd 14 13 pch_mac_CDNS_4618498380414 $T=10950 25305 0 0 $X=10170 $Y=24945
.ENDS
***************************************
.SUBCKT nch_CDNS_461849838041 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=1e-07 W=2e-07 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_CDNS_461849838040 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=1e-07 W=2e-07 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT rppolywo_CDNS_4618498380417 1 2
** N=3 EP=2 IP=0 FDC=1
X0 1 2 rppolywo l=8.534e-05 w=5e-07 $X=410 $Y=0 $D=215
.ENDS
***************************************
.SUBCKT ladder_R Rb Ra
** N=6 EP=2 IP=12 FDC=4
X0 Rb 5 rppolywo_CDNS_4618498380417 $T=8430 15120 0 0 $X=8230 $Y=14900
X1 4 5 rppolywo_CDNS_4618498380417 $T=8430 16550 0 0 $X=8230 $Y=16330
X2 4 6 rppolywo_CDNS_4618498380417 $T=8430 17990 0 0 $X=8230 $Y=17770
X3 Ra 6 rppolywo_CDNS_4618498380417 $T=8430 19430 0 0 $X=8230 $Y=19210
.ENDS
***************************************
.SUBCKT ladder_2R Rb Ra
** N=4 EP=2 IP=6 FDC=8
X0 Rb 4 ladder_R $T=-7360 -14095 0 0 $X=870 $Y=805
X1 4 Ra ladder_R $T=-7360 -8325 0 0 $X=870 $Y=6575
.ENDS
***************************************
.SUBCKT pch_CDNS_4618498380418 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=1e-07 W=2.5e-06 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4
** N=5 EP=4 IP=8 FDC=2
X0 2 1 3 pch_CDNS_461849838040 $T=0 0 0 0 $X=-780 $Y=-520
X1 2 4 1 pch_CDNS_4618498380418 $T=0 1445 0 0 $X=-780 $Y=925
.ENDS
***************************************
.SUBCKT nch_CDNS_4618498380421 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=1e-07 W=2.5e-06 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT nch_CDNS_4618498380420 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=1e-07 W=2e-07 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=11 FDC=4
X0 1 4 5 6 ICV_1 $T=0 0 0 0 $X=-780 $Y=-520
X1 2 7 3 nch_CDNS_4618498380421 $T=-1780 3945 0 180 $X=-2240 $Y=925
X2 2 3 8 nch_CDNS_4618498380420 $T=-1780 200 0 180 $X=-2240 $Y=-520
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=16 FDC=8
X0 3 2 1 7 8 9 5 6 ICV_2 $T=-2905 0 0 0 $X=-5145 $Y=-520
X1 4 2 3 7 10 11 9 8 ICV_2 $T=0 0 0 0 $X=-2240 $Y=-520
.ENDS
***************************************
.SUBCKT dac_real_res GND VREF B<1> B<2> B<6> B<3> B<5> B<7> B<0> B<4> VOUT
** N=34 EP=11 IP=97 FDC=132
M0 12 14 GND GND nch L=1e-07 W=2.5e-06 $X=7435 $Y=12240 $D=28
X1 29 28 ladder_R $T=8520 51635 1 0 $X=16750 $Y=31485
X2 30 29 ladder_R $T=8520 71125 1 0 $X=16750 $Y=50975
X3 31 30 ladder_R $T=8520 90615 1 0 $X=16750 $Y=70465
X4 32 31 ladder_R $T=102195 26395 1 0 $X=110425 $Y=6245
X5 33 32 ladder_R $T=102195 45875 1 0 $X=110425 $Y=25725
X6 34 33 ladder_R $T=102195 65355 1 0 $X=110425 $Y=45205
X7 VOUT 34 ladder_R $T=102195 84835 1 0 $X=110425 $Y=64685
X8 28 GND ladder_2R $T=15880 18050 1 0 $X=16750 $Y=6225
X9 28 12 ladder_2R $T=15880 18050 0 0 $X=16750 $Y=18855
X10 29 27 ladder_2R $T=15880 37540 0 0 $X=16750 $Y=38345
X11 30 26 ladder_2R $T=15880 57030 0 0 $X=16750 $Y=57835
X12 31 25 ladder_2R $T=15880 76520 0 0 $X=16750 $Y=77325
X13 32 23 ladder_2R $T=109555 12295 0 0 $X=110425 $Y=13100
X14 33 22 ladder_2R $T=109555 31775 0 0 $X=110425 $Y=32580
X15 34 21 ladder_2R $T=109555 51255 0 0 $X=110425 $Y=52060
X16 VOUT 24 ladder_2R $T=109555 70735 0 0 $X=110425 $Y=71540
X17 13 VREF B<7> 24 ICV_1 $T=5990 33700 0 270 $X=5470 $Y=33150
X18 GND 14 B<0> nch_CDNS_4618498380420 $T=6190 12240 0 90 $X=5470 $Y=11880
X19 15 GND 13 VREF B<6> 21 24 B<7> ICV_2 $T=5990 30795 0 270 $X=5470 $Y=30245
X20 16 GND 17 14 26 B<2> VREF B<1> 27 B<0> 12 ICV_3 $T=5990 13365 0 270 $X=5470 $Y=12815
X21 18 GND 19 16 23 B<4> VREF B<3> 25 B<2> 26 ICV_3 $T=5990 19175 0 270 $X=5470 $Y=18625
X22 15 GND 20 18 21 B<6> VREF B<5> 22 B<4> 23 ICV_3 $T=5990 24985 0 270 $X=5470 $Y=24435
.ENDS
***************************************
.SUBCKT pch_CDNS_461849838044 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 2 4 1 3 pch L=1e-07 W=2e-07 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_CDNS_461849838043 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=1e-07 W=2e-07 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_CDNS_461849838042 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=1e-07 W=2e-07 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT buffer OUT IN GND VDD
** N=5 EP=4 IP=14 FDC=4
X0 GND 5 IN nch_CDNS_461849838041 $T=830 800 0 90 $X=110 $Y=110
X1 GND OUT 5 nch_CDNS_461849838041 $T=1750 800 0 90 $X=1030 $Y=110
X2 VDD 5 IN pch_CDNS_461849838040 $T=630 2085 0 270 $X=110 $Y=1535
X3 VDD OUT 5 pch_CDNS_461849838040 $T=1550 2085 0 270 $X=1030 $Y=1535
.ENDS
***************************************
.SUBCKT SAR_system_3_u_sar_logic VIN GND VDD NQ B_Buf<0> B_Buf<1> B_Buf<2> B_Buf<3> B_Buf<4> B_Buf<5> B_Buf<6> B_Buf<7> VREF SoC EoC B<7> B<6> B<5> B<4> B<3>
+ B<2> B<1> B<0> COMP_OUT
** N=30 EP=24 IP=85 FDC=208
M0 2 7 VIN GND nch L=1e-07 W=2e-07 $X=40445 $Y=133500 $D=28
M1 2 6 VIN VDD pch L=1e-07 W=2e-07 $X=40445 $Y=134740 $D=62
X2 2 GND mimcap_2p0_sin lt=2.2065e-05 wt=2.2065e-05 $X=28215 $Y=123100 $D=151
X3 GND COMP_OUT VDD 2 30 comparator_rail2rail_input_external_current $T=65805 109620 0 0 $X=66720 $Y=110235
X4 GND NQ SoC nch_CDNS_461849838041 $T=11160 133640 0 180 $X=10700 $Y=132920
X5 GND 6 NQ nch_CDNS_461849838041 $T=14470 133640 0 180 $X=14010 $Y=132920
X6 GND 7 6 nch_CDNS_461849838041 $T=38480 133500 0 0 $X=37790 $Y=133140
X7 VDD 7 6 pch_CDNS_461849838040 $T=38480 134740 0 0 $X=37700 $Y=134220
X8 GND VREF B<6> B<5> B<1> B<4> B<2> B<0> B<7> B<3> 30 dac_real_res $T=19080 13900 0 0 $X=22630 $Y=20125
X9 8 NQ VDD SoC pch_CDNS_461849838044 $T=11060 134695 0 0 $X=10610 $Y=134335
X10 9 6 VDD NQ pch_CDNS_461849838044 $T=14370 134695 0 0 $X=13920 $Y=134335
X11 GND NQ 6 nch_CDNS_461849838043 $T=9860 133440 0 0 $X=9170 $Y=132920
X12 GND 6 EoC nch_CDNS_461849838043 $T=13125 133440 0 0 $X=12435 $Y=132920
X13 VDD 8 6 pch_CDNS_461849838042 $T=9860 134695 0 0 $X=9080 $Y=134335
X14 VDD 9 EoC pch_CDNS_461849838042 $T=13125 134695 0 0 $X=12345 $Y=134335
X15 B_Buf<0> B<7> GND VDD buffer $T=7175 25265 0 270 $X=7285 $Y=22725
X16 B_Buf<1> B<6> GND VDD buffer $T=7175 28860 0 270 $X=7285 $Y=26320
X17 B_Buf<2> B<5> GND VDD buffer $T=7175 32455 0 270 $X=7285 $Y=29915
X18 B_Buf<3> B<4> GND VDD buffer $T=7175 36050 0 270 $X=7285 $Y=33510
X19 B_Buf<4> B<3> GND VDD buffer $T=7175 39645 0 270 $X=7285 $Y=37105
X20 B_Buf<5> B<2> GND VDD buffer $T=7175 43240 0 270 $X=7285 $Y=40700
X21 B_Buf<6> B<1> GND VDD buffer $T=7175 46835 0 270 $X=7285 $Y=44295
X22 B_Buf<7> B<0> GND VDD buffer $T=7175 50430 0 270 $X=7285 $Y=47890
.ENDS
***************************************
