* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461414680674 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=2e-07 W=2e-06 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461414680676 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=1e-07 W=2e-06 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461414680671 1 2
** N=3 EP=2 IP=0 FDC=1
M0 2 2 1 1 pch L=1e-07 W=2e-06 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461414680670 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 pch L=5e-07 W=2e-06 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461414680679 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=1e-07 W=2.03e-06 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_4614146806711 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=1e-07 W=2e-06 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461414680678 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=2e-07 W=2e-06 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT comparator_rail2rail_input_external_current_small Gnd Vdd Out I_b I_t Ref In
** N=14 EP=7 IP=86 FDC=29
M0 3 In 2 Gnd nch L=5e-07 W=2e-06 $X=13390 $Y=4040 $D=28
M1 4 Ref 2 Gnd nch L=5e-07 W=2e-06 $X=14880 $Y=4040 $D=28
M2 6 I_b Gnd Gnd nch L=2e-07 W=1e-06 $X=16990 $Y=5165 $D=28
M3 Out 6 Gnd Gnd nch L=5e-07 W=1e-06 $X=17910 $Y=5165 $D=28
M4 Out 6 Vdd Vdd pch L=5e-07 W=2e-06 $X=17520 $Y=7470 $D=62
X5 Gnd 2 I_b nch_mac_CDNS_461414680674 $T=16990 1850 0 0 $X=16630 $Y=1490
X6 Gnd I_b I_b nch_mac_CDNS_461414680674 $T=18470 1845 0 0 $X=18110 $Y=1485
X7 Vdd 3 3 pch_mac_CDNS_461414680676 $T=4220 7470 0 0 $X=3440 $Y=7110
X8 Vdd 4 4 pch_mac_CDNS_461414680676 $T=13530 7470 0 0 $X=12750 $Y=7110
X9 Vdd 6 4 pch_mac_CDNS_461414680676 $T=14860 7470 0 0 $X=14080 $Y=7110
X10 Vdd 6 4 pch_mac_CDNS_461414680676 $T=16190 7470 0 0 $X=15410 $Y=7110
X11 Vdd 3 pch_mac_CDNS_461414680671 $T=5550 7470 0 0 $X=4770 $Y=6950
X12 Vdd 4 pch_mac_CDNS_461414680671 $T=12200 7470 0 0 $X=11420 $Y=6950
X13 Vdd 12 9 Ref pch_mac_CDNS_461414680670 $T=9095 4045 0 0 $X=8145 $Y=3525
X14 Vdd 12 10 In pch_mac_CDNS_461414680670 $T=11180 4045 0 0 $X=10230 $Y=3525
X15 Vdd 4 3 pch_mac_CDNS_461414680679 $T=6880 7440 0 0 $X=6100 $Y=7080
X16 Vdd 4 3 pch_mac_CDNS_461414680679 $T=8210 7440 0 0 $X=7430 $Y=7080
X17 Vdd 3 4 pch_mac_CDNS_461414680679 $T=9540 7440 0 0 $X=8760 $Y=7080
X18 Vdd 3 4 pch_mac_CDNS_461414680679 $T=10870 7440 0 0 $X=10090 $Y=7080
X19 Gnd 10 10 nch_mac_CDNS_4614146806711 $T=3355 2085 0 90 $X=995 $Y=1725
X20 Gnd 10 10 nch_mac_CDNS_4614146806711 $T=3355 3175 0 90 $X=995 $Y=2815
X21 Gnd 4 10 nch_mac_CDNS_4614146806711 $T=3355 4265 0 90 $X=995 $Y=3905
X22 Gnd 4 10 nch_mac_CDNS_4614146806711 $T=3355 5355 0 90 $X=995 $Y=4995
X23 Gnd 3 9 nch_mac_CDNS_4614146806711 $T=7290 2085 0 90 $X=4930 $Y=1725
X24 Gnd 3 9 nch_mac_CDNS_4614146806711 $T=7290 3175 0 90 $X=4930 $Y=2815
X25 Gnd 9 9 nch_mac_CDNS_4614146806711 $T=7290 4265 0 90 $X=4930 $Y=3905
X26 Gnd 9 9 nch_mac_CDNS_4614146806711 $T=7290 5355 0 90 $X=4930 $Y=4995
X27 Vdd I_t I_t pch_mac_CDNS_461414680678 $T=1360 7470 0 0 $X=580 $Y=7110
X28 Vdd 12 I_t pch_mac_CDNS_461414680678 $T=2790 7470 0 0 $X=2010 $Y=7110
.ENDS
***************************************
