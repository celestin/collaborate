* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461775247985 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=1e-06 W=2e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461775247987 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 4 1 3 nch L=5e-07 W=2e-06 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_4617752479810 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 2 4 1 3 pch L=5e-07 W=2e-06 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461775247980 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=2e-06 W=5e-06 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461775247982 1 2
** N=3 EP=2 IP=0 FDC=1
M0 2 2 1 1 pch L=1e-06 W=2e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_4617752479811 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=2e-06 W=2e-05 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461775247984 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=1e-06 W=2.03e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461775247983 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=1e-06 W=2e-05 $X=0 $Y=0 $D=28
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461775247989 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=2e-06 W=2e-05 $X=0 $Y=0 $D=62
.ENDS
***************************************
.SUBCKT comparator_rail2rail_input_external_current Gnd Out Vdd In Ref
** N=14 EP=5 IP=100 FDC=31
M0 Out 7 Gnd Gnd nch L=5e-07 W=1e-06 $X=31695 $Y=22735 $D=28
M1 Out 7 Vdd Vdd pch L=5e-07 W=2e-06 $X=33660 $Y=21735 $D=62
X2 8 11 rppolywo l=3.831e-05 w=8e-07 $X=4870 $Y=2205 $D=215
X3 Vdd 5 5 pch_mac_CDNS_461775247985 $T=14180 25305 0 0 $X=13400 $Y=24945
X4 Vdd 6 6 pch_mac_CDNS_461775247985 $T=29790 25305 0 0 $X=29010 $Y=24945
X5 Vdd 7 6 pch_mac_CDNS_461775247985 $T=32020 25305 0 0 $X=31240 $Y=24945
X6 Vdd 7 6 pch_mac_CDNS_461775247985 $T=34250 25305 0 0 $X=33470 $Y=24945
X7 4 5 Gnd In nch_mac_CDNS_461775247987 $T=29290 1960 0 0 $X=28930 $Y=1600
X8 4 6 Gnd Ref nch_mac_CDNS_461775247987 $T=31280 1960 0 0 $X=30920 $Y=1600
X9 12 9 Vdd In pch_mac_CDNS_4617752479810 $T=29335 18665 0 0 $X=28885 $Y=18145
X10 12 10 Vdd Ref pch_mac_CDNS_4617752479810 $T=31235 18665 0 0 $X=30785 $Y=18145
X11 Gnd 7 8 nch_mac_CDNS_461775247980 $T=29290 5860 0 0 $X=28930 $Y=5340
X12 Gnd 7 8 nch_mac_CDNS_461775247980 $T=29290 12195 0 0 $X=28930 $Y=11675
X13 Vdd 5 pch_mac_CDNS_461775247982 $T=16410 25305 0 0 $X=15630 $Y=24785
X14 Vdd 6 pch_mac_CDNS_461775247982 $T=27560 25305 0 0 $X=26780 $Y=24785
X15 Gnd 8 8 nch_mac_CDNS_4617752479811 $T=23310 1960 0 0 $X=22950 $Y=1600
X16 Gnd 4 8 nch_mac_CDNS_4617752479811 $T=26300 1960 0 0 $X=25940 $Y=1600
X17 Vdd 6 5 pch_mac_CDNS_461775247984 $T=18640 25005 0 0 $X=17860 $Y=24645
X18 Vdd 6 5 pch_mac_CDNS_461775247984 $T=20870 25005 0 0 $X=20090 $Y=24645
X19 Vdd 5 6 pch_mac_CDNS_461775247984 $T=23100 25005 0 0 $X=22320 $Y=24645
X20 Vdd 5 6 pch_mac_CDNS_461775247984 $T=25330 25005 0 0 $X=24550 $Y=24645
X21 Gnd 9 9 nch_mac_CDNS_461775247983 $T=7390 1955 0 0 $X=7030 $Y=1595
X22 Gnd 9 9 nch_mac_CDNS_461775247983 $T=9380 1955 0 0 $X=9020 $Y=1595
X23 Gnd 6 9 nch_mac_CDNS_461775247983 $T=11370 1955 0 0 $X=11010 $Y=1595
X24 Gnd 6 9 nch_mac_CDNS_461775247983 $T=13360 1955 0 0 $X=13000 $Y=1595
X25 Gnd 5 10 nch_mac_CDNS_461775247983 $T=15350 1955 0 0 $X=14990 $Y=1595
X26 Gnd 5 10 nch_mac_CDNS_461775247983 $T=17340 1955 0 0 $X=16980 $Y=1595
X27 Gnd 10 10 nch_mac_CDNS_461775247983 $T=19330 1955 0 0 $X=18970 $Y=1595
X28 Gnd 10 10 nch_mac_CDNS_461775247983 $T=21320 1955 0 0 $X=20960 $Y=1595
X29 Vdd 11 11 pch_mac_CDNS_461775247989 $T=7720 25305 0 0 $X=6940 $Y=24945
X30 Vdd 12 11 pch_mac_CDNS_461775247989 $T=10950 25305 0 0 $X=10170 $Y=24945
.ENDS
***************************************
