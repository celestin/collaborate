* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_2p0_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_4619242438510
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_4619242438512
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_4619242438515
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461924243855
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461924243857
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_4619242438516
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_461924243859
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_mac_CDNS_461924243858
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pch_mac_CDNS_4619242438514
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT comparator_rail2rail_input_external_current Gnd Out Vdd In Ref
** N=14 EP=5 IP=100 FDC=31
M0 Out 9 Gnd Gnd nch L=5e-07 W=1e-06 AD=2.3e-13 AS=2.3e-13 PD=2.46e-06 PS=2.46e-06 NRD=0.23 NRS=0.23 sa=2.3e-07 sb=2.3e-07 sca=1.77318 scb=0.000164701 scc=8.24936e-08 $X=31695 $Y=22735 $D=28
M1 7 In 6 Gnd nch L=5e-07 W=2e-06 AD=4.6e-13 AS=4.6e-13 PD=4.46e-06 PS=4.46e-06 NRD=0.115 NRS=0.115 sa=2.3e-07 sb=2.3e-07 sca=0.12987 scb=4.8892e-22 scc=4.69641e-44 $X=29290 $Y=1960 $D=28
M2 8 Ref 6 Gnd nch L=5e-07 W=2e-06 AD=4.6e-13 AS=4.6e-13 PD=4.46e-06 PS=4.46e-06 NRD=0.115 NRS=0.115 sa=2.3e-07 sb=2.3e-07 sca=0.12987 scb=4.8892e-22 scc=4.69641e-44 $X=31280 $Y=1960 $D=28
M3 9 10 Gnd Gnd nch L=2e-06 W=5e-06 AD=1.15e-12 AS=1.15e-12 PD=1.046e-05 PS=1.046e-05 NRD=0.046 NRS=0.046 sa=2.3e-07 sb=2.3e-07 sca=0.0971429 scb=1.37713e-22 scc=1.31505e-44 $X=29290 $Y=5860 $D=28
M4 9 10 Gnd Gnd nch L=2e-06 W=5e-06 AD=1.15e-12 AS=1.15e-12 PD=1.046e-05 PS=1.046e-05 NRD=0.046 NRS=0.046 sa=2.3e-07 sb=2.3e-07 sca=0.205143 scb=1.0062e-07 scc=1.80543e-13 $X=29290 $Y=12195 $D=28
M5 10 10 Gnd Gnd nch L=2e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.0832869 scb=7.88215e-15 scc=2.0842e-27 $X=23310 $Y=1960 $D=28
M6 6 10 Gnd Gnd nch L=2e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.156674 scb=1.20337e-05 scc=1.60631e-08 $X=26300 $Y=1960 $D=28
M7 11 11 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.0884794 scb=4.11866e-16 scc=5.1705e-30 $X=7390 $Y=1955 $D=28
M8 11 11 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.0884794 scb=4.11866e-16 scc=5.1705e-30 $X=9380 $Y=1955 $D=28
M9 8 11 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.0884794 scb=4.11866e-16 scc=5.1705e-30 $X=11370 $Y=1955 $D=28
M10 8 11 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.0884794 scb=4.11866e-16 scc=5.1705e-30 $X=13360 $Y=1955 $D=28
M11 7 12 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.0884794 scb=4.11866e-16 scc=5.1705e-30 $X=15350 $Y=1955 $D=28
M12 7 12 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.0892786 scb=3.81618e-15 scc=9.09477e-28 $X=17340 $Y=1955 $D=28
M13 12 12 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.0901444 scb=7.50419e-15 scc=1.88914e-27 $X=19330 $Y=1955 $D=28
M14 12 12 Gnd Gnd nch L=1e-06 W=2e-05 AD=4.6e-12 AS=4.6e-12 PD=4.046e-05 PS=4.046e-05 NRD=0.0115 NRS=0.0115 sa=2.3e-07 sb=2.3e-07 sca=0.0901444 scb=7.50419e-15 scc=1.88914e-27 $X=21320 $Y=1955 $D=28
M15 Out 9 Vdd Vdd pch L=5e-07 W=2e-06 AD=4.6e-13 AS=6.4e-13 PD=4.46e-06 PS=4.64e-06 NRD=0.115 NRS=0.16 sa=5.6e-07 sb=2.3e-07 sca=7.43579 scb=0.00482332 scc=0.000171928 $X=33660 $Y=21735 $D=62
M16 7 7 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.516267 scb=0.00035457 scc=1.65744e-05 $X=14180 $Y=25305 $D=62
M17 8 8 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.517394 scb=0.00035457 scc=1.65744e-05 $X=29790 $Y=25305 $D=62
M18 9 8 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.584328 scb=0.00035457 scc=1.65744e-05 $X=32020 $Y=25305 $D=62
M19 9 8 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=2.0155 scb=0.000965487 scc=1.96597e-05 $X=34250 $Y=25305 $D=62
M20 11 In 14 Vdd pch L=5e-07 W=2e-06 AD=4.6e-13 AS=4.6e-13 PD=4.46e-06 PS=4.46e-06 NRD=0.115 NRS=0.115 sa=2.3e-07 sb=2.3e-07 sca=6.53892 scb=0.00475197 scc=0.000171914 $X=29335 $Y=18665 $D=62
M21 12 Ref 14 Vdd pch L=5e-07 W=2e-06 AD=4.6e-13 AS=4.6e-13 PD=4.46e-06 PS=4.46e-06 NRD=0.115 NRS=0.115 sa=2.3e-07 sb=2.3e-07 sca=4.97027 scb=0.00356126 scc=0.000165745 $X=31235 $Y=18665 $D=62
M22 7 7 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.516267 scb=0.00035457 scc=1.65744e-05 $X=16410 $Y=25305 $D=62
M23 8 8 Vdd Vdd pch L=1e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.516267 scb=0.00035457 scc=1.65744e-05 $X=27560 $Y=25305 $D=62
M24 8 7 Vdd Vdd pch L=1e-06 W=2.03e-05 AD=4.669e-12 AS=6.496e-12 PD=4.106e-05 PS=4.124e-05 NRD=0.01133 NRS=0.0157635 sa=5.6e-07 sb=2.3e-07 sca=0.512401 scb=0.000349472 scc=1.63295e-05 $X=18640 $Y=25005 $D=62
M25 8 7 Vdd Vdd pch L=1e-06 W=2.03e-05 AD=4.669e-12 AS=6.496e-12 PD=4.106e-05 PS=4.124e-05 NRD=0.01133 NRS=0.0157635 sa=5.6e-07 sb=2.3e-07 sca=0.509893 scb=0.00034933 scc=1.63295e-05 $X=20870 $Y=25005 $D=62
M26 7 8 Vdd Vdd pch L=1e-06 W=2.03e-05 AD=4.669e-12 AS=6.496e-12 PD=4.106e-05 PS=4.124e-05 NRD=0.01133 NRS=0.0157635 sa=5.6e-07 sb=2.3e-07 sca=0.509962 scb=0.00034933 scc=1.63295e-05 $X=23100 $Y=25005 $D=62
M27 7 8 Vdd Vdd pch L=1e-06 W=2.03e-05 AD=4.669e-12 AS=6.496e-12 PD=4.106e-05 PS=4.124e-05 NRD=0.01133 NRS=0.0157635 sa=5.6e-07 sb=2.3e-07 sca=0.515602 scb=0.000351738 scc=1.63416e-05 $X=25330 $Y=25005 $D=62
M28 13 13 Vdd Vdd pch L=2e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.939341 scb=0.000372598 scc=1.65779e-05 $X=7720 $Y=25305 $D=62
M29 14 13 Vdd Vdd pch L=2e-06 W=2e-05 AD=4.6e-12 AS=6.4e-12 PD=4.046e-05 PS=4.064e-05 NRD=0.0115 NRS=0.016 sa=5.6e-07 sb=2.3e-07 sca=0.519665 scb=0.00035457 scc=1.65744e-05 $X=10950 $Y=25305 $D=62
X30 10 13 rppolywo l=3.831e-05 w=8e-07 $X=4870 $Y=2205 $D=215
.ENDS
***************************************
.SUBCKT nch_CDNS_461924243851
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pch_CDNS_461924243850
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT rppolywo_CDNS_4619242438517 1 2
** N=3 EP=2 IP=0 FDC=1
X0 1 2 rppolywo l=8.534e-05 w=5e-07 $X=410 $Y=0 $D=215
.ENDS
***************************************
.SUBCKT ladder_R Rb Ra
** N=6 EP=2 IP=12 FDC=4
X0 Rb 5 rppolywo_CDNS_4619242438517 $T=8430 15120 0 0 $X=8230 $Y=14900
X1 4 5 rppolywo_CDNS_4619242438517 $T=8430 16550 0 0 $X=8230 $Y=16330
X2 4 6 rppolywo_CDNS_4619242438517 $T=8430 17990 0 0 $X=8230 $Y=17770
X3 Ra 6 rppolywo_CDNS_4619242438517 $T=8430 19430 0 0 $X=8230 $Y=19210
.ENDS
***************************************
.SUBCKT ladder_2R Rb Ra
** N=4 EP=2 IP=6 FDC=8
X0 Rb 4 ladder_R $T=-7360 -14095 0 0 $X=870 $Y=805
X1 4 Ra ladder_R $T=-7360 -8325 0 0 $X=870 $Y=6575
.ENDS
***************************************
.SUBCKT pch_CDNS_4619242438518
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_1
** N=5 EP=0 IP=7 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_CDNS_4619242438521
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_CDNS_4619242438520
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_2
** N=8 EP=0 IP=11 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_3
** N=11 EP=0 IP=16 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT dac_real_res GND VREF B<1> B<2> B<6> B<3> B<5> B<7> B<0> B<4> VOUT
** N=34 EP=11 IP=97 FDC=132
M0 12 14 GND GND nch L=1e-07 W=2.5e-06 AD=5.75e-13 AS=8e-13 PD=5.46e-06 PS=5.64e-06 NRD=0.092 NRS=0.128 sa=5.6e-07 sb=2.3e-07 sca=3.75388 scb=0.00282635 scc=1.6483e-05 $X=7435 $Y=12240 $D=28
M1 14 B<0> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=3.77747 scb=0.00282635 scc=1.6483e-05 $X=5990 $Y=12240 $D=28
M2 24 13 GND GND nch L=1e-07 W=2.5e-06 AD=5.75e-13 AS=5.75e-13 PD=5.46e-06 PS=5.46e-06 NRD=0.092 NRS=0.092 sa=2.3e-07 sb=2.3e-07 sca=4.62375 scb=0.00285625 scc=1.64839e-05 $X=7435 $Y=32575 $D=28
M3 13 B<7> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=4.64734 scb=0.00285625 scc=1.64839e-05 $X=5990 $Y=32575 $D=28
M4 26 16 GND GND nch L=1e-07 W=2.5e-06 AD=5.75e-13 AS=5.75e-13 PD=5.46e-06 PS=5.46e-06 NRD=0.092 NRS=0.092 sa=2.3e-07 sb=2.3e-07 sca=4.62375 scb=0.00285625 scc=1.64839e-05 $X=7435 $Y=18050 $D=28
M5 16 B<2> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=4.64734 scb=0.00285625 scc=1.64839e-05 $X=5990 $Y=18050 $D=28
M6 27 17 GND GND nch L=1e-07 W=2.5e-06 AD=5.75e-13 AS=5.75e-13 PD=5.46e-06 PS=5.46e-06 NRD=0.092 NRS=0.092 sa=2.3e-07 sb=2.3e-07 sca=4.62375 scb=0.00285625 scc=1.64839e-05 $X=7435 $Y=15145 $D=28
M7 17 B<1> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=4.64734 scb=0.00285625 scc=1.64839e-05 $X=5990 $Y=15145 $D=28
M8 23 18 GND GND nch L=1e-07 W=2.5e-06 AD=5.75e-13 AS=5.75e-13 PD=5.46e-06 PS=5.46e-06 NRD=0.092 NRS=0.092 sa=2.3e-07 sb=2.3e-07 sca=4.62375 scb=0.00285625 scc=1.64839e-05 $X=7435 $Y=23860 $D=28
M9 18 B<4> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=4.64734 scb=0.00285625 scc=1.64839e-05 $X=5990 $Y=23860 $D=28
M10 25 19 GND GND nch L=1e-07 W=2.5e-06 AD=5.75e-13 AS=5.75e-13 PD=5.46e-06 PS=5.46e-06 NRD=0.092 NRS=0.092 sa=2.3e-07 sb=2.3e-07 sca=4.62375 scb=0.00285625 scc=1.64839e-05 $X=7435 $Y=20955 $D=28
M11 19 B<3> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=4.64734 scb=0.00285625 scc=1.64839e-05 $X=5990 $Y=20955 $D=28
M12 21 15 GND GND nch L=1e-07 W=2.5e-06 AD=5.75e-13 AS=5.75e-13 PD=5.46e-06 PS=5.46e-06 NRD=0.092 NRS=0.092 sa=2.3e-07 sb=2.3e-07 sca=4.62375 scb=0.00285625 scc=1.64839e-05 $X=7435 $Y=29670 $D=28
M13 15 B<6> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=4.64734 scb=0.00285625 scc=1.64839e-05 $X=5990 $Y=29670 $D=28
M14 22 20 GND GND nch L=1e-07 W=2.5e-06 AD=5.75e-13 AS=5.75e-13 PD=5.46e-06 PS=5.46e-06 NRD=0.092 NRS=0.092 sa=2.3e-07 sb=2.3e-07 sca=4.62375 scb=0.00285625 scc=1.64839e-05 $X=7435 $Y=26765 $D=28
M15 20 B<5> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=4.64734 scb=0.00285625 scc=1.64839e-05 $X=5990 $Y=26765 $D=28
M16 VREF B<7> 13 VREF pch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=16.3803 scb=0.0174961 scc=0.0008282 $X=5990 $Y=33600 $D=62
M17 VREF 13 24 VREF pch L=1e-07 W=2.5e-06 AD=8e-13 AS=5.75e-13 PD=5.64e-06 PS=5.46e-06 NRD=0.128 NRS=0.092 sa=2.3e-07 sb=5.6e-07 sca=7.31261 scb=0.00508468 scc=9.21987e-05 $X=7435 $Y=33600 $D=62
M18 VREF B<6> 15 VREF pch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=16.3803 scb=0.0174961 scc=0.0008282 $X=5990 $Y=30695 $D=62
M19 VREF 15 21 VREF pch L=1e-07 W=2.5e-06 AD=8e-13 AS=5.75e-13 PD=5.64e-06 PS=5.46e-06 NRD=0.128 NRS=0.092 sa=2.3e-07 sb=5.6e-07 sca=7.31261 scb=0.00508468 scc=9.21987e-05 $X=7435 $Y=30695 $D=62
M20 VREF B<1> 17 VREF pch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=16.3803 scb=0.0174961 scc=0.0008282 $X=5990 $Y=16170 $D=62
M21 VREF 17 27 VREF pch L=1e-07 W=2.5e-06 AD=8e-13 AS=5.75e-13 PD=5.64e-06 PS=5.46e-06 NRD=0.128 NRS=0.092 sa=2.3e-07 sb=5.6e-07 sca=7.31261 scb=0.00508468 scc=9.21987e-05 $X=7435 $Y=16170 $D=62
M22 VREF B<0> 14 VREF pch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=16.3803 scb=0.0174961 scc=0.0008282 $X=5990 $Y=13265 $D=62
M23 VREF 14 12 VREF pch L=1e-07 W=2.5e-06 AD=8e-13 AS=5.75e-13 PD=5.64e-06 PS=5.46e-06 NRD=0.128 NRS=0.092 sa=2.3e-07 sb=5.6e-07 sca=7.31261 scb=0.00508468 scc=9.21987e-05 $X=7435 $Y=13265 $D=62
M24 VREF B<3> 19 VREF pch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=16.3803 scb=0.0174961 scc=0.0008282 $X=5990 $Y=21980 $D=62
M25 VREF 19 25 VREF pch L=1e-07 W=2.5e-06 AD=8e-13 AS=5.75e-13 PD=5.64e-06 PS=5.46e-06 NRD=0.128 NRS=0.092 sa=2.3e-07 sb=5.6e-07 sca=7.31261 scb=0.00508468 scc=9.21987e-05 $X=7435 $Y=21980 $D=62
M26 VREF B<2> 16 VREF pch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=16.3803 scb=0.0174961 scc=0.0008282 $X=5990 $Y=19075 $D=62
M27 VREF 16 26 VREF pch L=1e-07 W=2.5e-06 AD=8e-13 AS=5.75e-13 PD=5.64e-06 PS=5.46e-06 NRD=0.128 NRS=0.092 sa=2.3e-07 sb=5.6e-07 sca=7.31261 scb=0.00508468 scc=9.21987e-05 $X=7435 $Y=19075 $D=62
M28 VREF B<5> 20 VREF pch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=16.3803 scb=0.0174961 scc=0.0008282 $X=5990 $Y=27790 $D=62
M29 VREF 20 22 VREF pch L=1e-07 W=2.5e-06 AD=8e-13 AS=5.75e-13 PD=5.64e-06 PS=5.46e-06 NRD=0.128 NRS=0.092 sa=2.3e-07 sb=5.6e-07 sca=7.31261 scb=0.00508468 scc=9.21987e-05 $X=7435 $Y=27790 $D=62
M30 VREF B<4> 18 VREF pch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=16.3803 scb=0.0174961 scc=0.0008282 $X=5990 $Y=24885 $D=62
M31 VREF 18 23 VREF pch L=1e-07 W=2.5e-06 AD=8e-13 AS=5.75e-13 PD=5.64e-06 PS=5.46e-06 NRD=0.128 NRS=0.092 sa=2.3e-07 sb=5.6e-07 sca=7.31261 scb=0.00508468 scc=9.21987e-05 $X=7435 $Y=24885 $D=62
X32 29 28 ladder_R $T=8520 51635 1 0 $X=16750 $Y=31485
X33 30 29 ladder_R $T=8520 71125 1 0 $X=16750 $Y=50975
X34 31 30 ladder_R $T=8520 90615 1 0 $X=16750 $Y=70465
X35 32 31 ladder_R $T=102195 26395 1 0 $X=110425 $Y=6245
X36 33 32 ladder_R $T=102195 45875 1 0 $X=110425 $Y=25725
X37 34 33 ladder_R $T=102195 65355 1 0 $X=110425 $Y=45205
X38 VOUT 34 ladder_R $T=102195 84835 1 0 $X=110425 $Y=64685
X39 28 GND ladder_2R $T=15880 18050 1 0 $X=16750 $Y=6225
X40 28 12 ladder_2R $T=15880 18050 0 0 $X=16750 $Y=18855
X41 29 27 ladder_2R $T=15880 37540 0 0 $X=16750 $Y=38345
X42 30 26 ladder_2R $T=15880 57030 0 0 $X=16750 $Y=57835
X43 31 25 ladder_2R $T=15880 76520 0 0 $X=16750 $Y=77325
X44 32 23 ladder_2R $T=109555 12295 0 0 $X=110425 $Y=13100
X45 33 22 ladder_2R $T=109555 31775 0 0 $X=110425 $Y=32580
X46 34 21 ladder_2R $T=109555 51255 0 0 $X=110425 $Y=52060
X47 VOUT 24 ladder_2R $T=109555 70735 0 0 $X=110425 $Y=71540
.ENDS
***************************************
.SUBCKT pch_CDNS_461924243854
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nch_CDNS_461924243853
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pch_CDNS_461924243852
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT buffer OUT IN VDD 5
** N=5 EP=4 IP=12 FDC=2
*.SEEDPROM
M0 VDD IN 5 VDD pch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=7.53827 scb=0.00345363 scc=1.14707e-05 $X=630 $Y=1985 $D=62
M1 VDD 5 OUT VDD pch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=8.26369 scb=0.0045196 scc=2.02638e-05 $X=1550 $Y=1985 $D=62
.ENDS
***************************************
.SUBCKT SAR_system_3_u_sar_logic VIN GND VDD NQ B_Buf<0> B_Buf<1> B_Buf<2> B_Buf<3> B_Buf<4> B_Buf<5> B_Buf<6> B_Buf<7> VREF SoC EoC B<7> B<6> B<5> B<4> B<3>
+ B<2> B<1> B<0> COMP_OUT
** N=38 EP=24 IP=92 FDC=208
M0 2 7 VIN GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=1.31249 scb=0.000105525 scc=1.60374e-08 $X=40445 $Y=133500 $D=28
M1 GND SoC NQ GND nch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=1.50381 scb=0.000187353 scc=5.44306e-08 $X=11060 $Y=133440 $D=28
M2 GND NQ 6 GND nch L=1e-07 W=2e-07 AD=6.4e-14 AS=4.6e-14 PD=1.04e-06 PS=8.6e-07 NRD=1.6 NRS=1.15 sa=2.3e-07 sb=5.6e-07 sca=1.50381 scb=0.000187353 scc=5.44306e-08 $X=14370 $Y=133440 $D=28
M3 7 6 GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=1.31249 scb=0.000105525 scc=1.60374e-08 $X=38480 $Y=133500 $D=28
M4 NQ 6 GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=1.50381 scb=0.000187353 scc=5.44306e-08 $X=9860 $Y=133440 $D=28
M5 6 EoC GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=1.50381 scb=0.000187353 scc=5.44306e-08 $X=13125 $Y=133440 $D=28
M6 31 B<7> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.7055 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=24435 $D=28
M7 B_Buf<0> 31 GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.7361 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=23515 $D=28
M8 32 B<6> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=28030 $D=28
M9 B_Buf<1> 32 GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=27110 $D=28
M10 33 B<5> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=31625 $D=28
M11 B_Buf<2> 33 GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=30705 $D=28
M12 34 B<4> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=35220 $D=28
M13 B_Buf<3> 34 GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=34300 $D=28
M14 35 B<3> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=38815 $D=28
M15 B_Buf<4> 35 GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=37895 $D=28
M16 36 B<2> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=42410 $D=28
M17 B_Buf<5> 36 GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=41490 $D=28
M18 37 B<1> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=46005 $D=28
M19 B_Buf<6> 37 GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=45085 $D=28
M20 38 B<0> GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=49600 $D=28
M21 B_Buf<7> 38 GND GND nch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=2.69263 scb=0.00124095 scc=2.66868e-06 $X=7975 $Y=48680 $D=28
M22 2 6 VIN VDD pch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=22.6484 scb=0.0276843 scc=0.0016046 $X=40445 $Y=134740 $D=62
M23 7 6 VDD VDD pch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=23.2105 scb=0.0278722 scc=0.00160466 $X=38480 $Y=134740 $D=62
M24 NQ SoC 8 VDD pch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=9.51618 scb=0.00922803 scc=0.000214172 $X=11060 $Y=134695 $D=62
M25 6 NQ 9 VDD pch L=1e-07 W=2e-07 AD=4.6e-14 AS=4.6e-14 PD=8.6e-07 PS=8.6e-07 NRD=1.15 NRS=1.15 sa=2.3e-07 sb=2.3e-07 sca=9.94725 scb=0.00923357 scc=0.000214172 $X=14370 $Y=134695 $D=62
M26 8 6 VDD VDD pch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=10.4016 scb=0.0093015 scc=0.000214178 $X=9860 $Y=134695 $D=62
M27 9 EoC VDD VDD pch L=1e-07 W=2e-07 AD=4.6e-14 AS=6.4e-14 PD=8.6e-07 PS=1.04e-06 NRD=1.15 NRS=1.6 sa=5.6e-07 sb=2.3e-07 sca=9.47027 scb=0.00922803 scc=0.000214172 $X=13125 $Y=134695 $D=62
X28 2 GND mimcap_2p0_sin lt=2.2065e-05 wt=2.2065e-05 $X=28215 $Y=123100 $D=151
X29 GND COMP_OUT VDD 2 30 comparator_rail2rail_input_external_current $T=65805 109620 0 0 $X=66720 $Y=110235
X34 GND VREF B<6> B<5> B<1> B<4> B<2> B<0> B<7> B<3> 30 dac_real_res $T=19080 13900 0 0 $X=22630 $Y=20125
X41 B_Buf<0> B<7> VDD 31 buffer $T=7175 25265 0 270 $X=7285 $Y=22725
X42 B_Buf<1> B<6> VDD 32 buffer $T=7175 28860 0 270 $X=7285 $Y=26320
X43 B_Buf<2> B<5> VDD 33 buffer $T=7175 32455 0 270 $X=7285 $Y=29915
X44 B_Buf<3> B<4> VDD 34 buffer $T=7175 36050 0 270 $X=7285 $Y=33510
X45 B_Buf<4> B<3> VDD 35 buffer $T=7175 39645 0 270 $X=7285 $Y=37105
X46 B_Buf<5> B<2> VDD 36 buffer $T=7175 43240 0 270 $X=7285 $Y=40700
X47 B_Buf<6> B<1> VDD 37 buffer $T=7175 46835 0 270 $X=7285 $Y=44295
X48 B_Buf<7> B<0> VDD 38 buffer $T=7175 50430 0 270 $X=7285 $Y=47890
.ENDS
***************************************
